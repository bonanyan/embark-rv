
module embarkrv (
    ports
);
    
endmodule